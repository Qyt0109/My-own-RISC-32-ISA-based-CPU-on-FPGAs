`include "global_constant.vh"

module RISC32_CPU (
    
);

endmodule //RISC32_CPU


